`timescale 1 ns / 100 ps
module lcd_ram(
        output reg [7:0] rom_q,
        input wire [8:0] rom_addr
);
	always @ (*)
		case(rom_addr)
            9'd0 : rom_q=8'hf8;
            9'd1 : rom_q=8'h0;
            9'd2 : rom_q=8'hf8;
            9'd3 : rom_q=8'h0;
            9'd4 : rom_q=8'hf8;
            9'd5 : rom_q=8'h0;
            9'd6 : rom_q=8'hf8;
            9'd7 : rom_q=8'h0;
            9'd8 : rom_q=8'hf8;
            9'd9 : rom_q=8'h0;
            9'd10 : rom_q=8'hf8;
            9'd11 : rom_q=8'h0;
            9'd12 : rom_q=8'hf8;
            9'd13 : rom_q=8'h0;
            9'd14 : rom_q=8'hf8;
            9'd15 : rom_q=8'h0;
            9'd16 : rom_q=8'hf8;
            9'd17 : rom_q=8'h0;
            9'd18 : rom_q=8'hf8;
            9'd19 : rom_q=8'h0;
            9'd20 : rom_q=8'hf8;
            9'd21 : rom_q=8'h0;
            9'd22 : rom_q=8'hf8;
            9'd23 : rom_q=8'h0;
            9'd24 : rom_q=8'hf8;
            9'd25 : rom_q=8'h0;
            9'd26 : rom_q=8'hf8;
            9'd27 : rom_q=8'h0;
            9'd28 : rom_q=8'hf8;
            9'd29 : rom_q=8'h0;
            9'd30 : rom_q=8'hf8;
            9'd31 : rom_q=8'h0;
            9'd32 : rom_q=8'hf8;
            9'd33 : rom_q=8'h0;
            9'd34 : rom_q=8'hf8;
            9'd35 : rom_q=8'h0;
            9'd36 : rom_q=8'hf8;
            9'd37 : rom_q=8'h0;
            9'd38 : rom_q=8'hf8;
            9'd39 : rom_q=8'h0;
            9'd40 : rom_q=8'hf8;
            9'd41 : rom_q=8'h0;
            9'd42 : rom_q=8'hf8;
            9'd43 : rom_q=8'h0;
            9'd44 : rom_q=8'hf8;
            9'd45 : rom_q=8'h0;
            9'd46 : rom_q=8'hf8;
            9'd47 : rom_q=8'h0;
            9'd48 : rom_q=8'hf8;
            9'd49 : rom_q=8'h0;
            9'd50 : rom_q=8'hf8;
            9'd51 : rom_q=8'h0;
            9'd52 : rom_q=8'hf8;
            9'd53 : rom_q=8'h0;
            9'd54 : rom_q=8'hf8;
            9'd55 : rom_q=8'h0;
            9'd56 : rom_q=8'hf8;
            9'd57 : rom_q=8'h0;
            9'd58 : rom_q=8'hf8;
            9'd59 : rom_q=8'h0;
            9'd60 : rom_q=8'hf8;
            9'd61 : rom_q=8'h0;
            9'd62 : rom_q=8'hf8;
            9'd63 : rom_q=8'h0;
            9'd64 : rom_q=8'hf8;
            9'd65 : rom_q=8'h0;
            9'd66 : rom_q=8'hf8;
            9'd67 : rom_q=8'h0;
            9'd68 : rom_q=8'hf8;
            9'd69 : rom_q=8'h0;
            9'd70 : rom_q=8'hf8;
            9'd71 : rom_q=8'h0;
            9'd72 : rom_q=8'hf8;
            9'd73 : rom_q=8'h0;
            9'd74 : rom_q=8'hf8;
            9'd75 : rom_q=8'h0;
            9'd76 : rom_q=8'hf8;
            9'd77 : rom_q=8'h0;
            9'd78 : rom_q=8'hf8;
            9'd79 : rom_q=8'h0;
            9'd80 : rom_q=8'hf8;
            9'd81 : rom_q=8'h0;
            9'd82 : rom_q=8'hf8;
            9'd83 : rom_q=8'h0;
            9'd84 : rom_q=8'hf8;
            9'd85 : rom_q=8'h0;
            9'd86 : rom_q=8'hf8;
            9'd87 : rom_q=8'h0;
            9'd88 : rom_q=8'hf8;
            9'd89 : rom_q=8'h0;
            9'd90 : rom_q=8'hf8;
            9'd91 : rom_q=8'h0;
            9'd92 : rom_q=8'hf8;
            9'd93 : rom_q=8'h0;
            9'd94 : rom_q=8'hf8;
            9'd95 : rom_q=8'h0;
            9'd96 : rom_q=8'hf8;
            9'd97 : rom_q=8'h0;
            9'd98 : rom_q=8'hf8;
            9'd99 : rom_q=8'h0;
            9'd100 : rom_q=8'hf8;
            9'd101 : rom_q=8'h0;
            9'd102 : rom_q=8'hf8;
            9'd103 : rom_q=8'h0;
            9'd104 : rom_q=8'hf8;
            9'd105 : rom_q=8'h0;
            9'd106 : rom_q=8'hf8;
            9'd107 : rom_q=8'h0;
            9'd108 : rom_q=8'hf8;
            9'd109 : rom_q=8'h0;
            9'd110 : rom_q=8'hf8;
            9'd111 : rom_q=8'h0;
            9'd112 : rom_q=8'hf8;
            9'd113 : rom_q=8'h0;
            9'd114 : rom_q=8'hf8;
            9'd115 : rom_q=8'h0;
            9'd116 : rom_q=8'hf8;
            9'd117 : rom_q=8'h0;
            9'd118 : rom_q=8'hf8;
            9'd119 : rom_q=8'h0;
            9'd120 : rom_q=8'hf8;
            9'd121 : rom_q=8'h0;
            9'd122 : rom_q=8'hf8;
            9'd123 : rom_q=8'h0;
            9'd124 : rom_q=8'hf8;
            9'd125 : rom_q=8'h0;
            9'd126 : rom_q=8'hf8;
            9'd127 : rom_q=8'h0;
            9'd128 : rom_q=8'hf8;
            9'd129 : rom_q=8'h0;
            9'd130 : rom_q=8'hf8;
            9'd131 : rom_q=8'h0;
            9'd132 : rom_q=8'hf8;
            9'd133 : rom_q=8'h0;
            9'd134 : rom_q=8'hf8;
            9'd135 : rom_q=8'h0;
            9'd136 : rom_q=8'hf8;
            9'd137 : rom_q=8'h0;
            9'd138 : rom_q=8'hf8;
            9'd139 : rom_q=8'h0;
            9'd140 : rom_q=8'hf8;
            9'd141 : rom_q=8'h0;
            9'd142 : rom_q=8'hf8;
            9'd143 : rom_q=8'h0;
            9'd144 : rom_q=8'hf8;
            9'd145 : rom_q=8'h0;
            9'd146 : rom_q=8'hf8;
            9'd147 : rom_q=8'h0;
            9'd148 : rom_q=8'hf8;
            9'd149 : rom_q=8'h0;
            9'd150 : rom_q=8'hf8;
            9'd151 : rom_q=8'h0;
            9'd152 : rom_q=8'hf8;
            9'd153 : rom_q=8'h0;
            9'd154 : rom_q=8'hf8;
            9'd155 : rom_q=8'h0;
            9'd156 : rom_q=8'hf8;
            9'd157 : rom_q=8'h0;
            9'd158 : rom_q=8'hf8;
            9'd159 : rom_q=8'h0;
            9'd160 : rom_q=8'hf8;
            9'd161 : rom_q=8'h0;
            9'd162 : rom_q=8'hf8;
            9'd163 : rom_q=8'h0;
            9'd164 : rom_q=8'hf8;
            9'd165 : rom_q=8'h0;
            9'd166 : rom_q=8'hf8;
            9'd167 : rom_q=8'h0;
            9'd168 : rom_q=8'hf8;
            9'd169 : rom_q=8'h0;
            9'd170 : rom_q=8'hf8;
            9'd171 : rom_q=8'h0;
            9'd172 : rom_q=8'hf8;
            9'd173 : rom_q=8'h0;
            9'd174 : rom_q=8'hf8;
            9'd175 : rom_q=8'h0;
            9'd176 : rom_q=8'hf8;
            9'd177 : rom_q=8'h0;
            9'd178 : rom_q=8'hf8;
            9'd179 : rom_q=8'h0;
            9'd180 : rom_q=8'hf8;
            9'd181 : rom_q=8'h0;
            9'd182 : rom_q=8'hf8;
            9'd183 : rom_q=8'h0;
            9'd184 : rom_q=8'hf8;
            9'd185 : rom_q=8'h0;
            9'd186 : rom_q=8'hf8;
            9'd187 : rom_q=8'h0;
            9'd188 : rom_q=8'hf8;
            9'd189 : rom_q=8'h0;
            9'd190 : rom_q=8'hf8;
            9'd191 : rom_q=8'h0;
            9'd192 : rom_q=8'hf8;
            9'd193 : rom_q=8'h0;
            9'd194 : rom_q=8'hf8;
            9'd195 : rom_q=8'h0;
            9'd196 : rom_q=8'hf8;
            9'd197 : rom_q=8'h0;
            9'd198 : rom_q=8'hf8;
            9'd199 : rom_q=8'h0;
            9'd200 : rom_q=8'hf8;
            9'd201 : rom_q=8'h0;
            9'd202 : rom_q=8'hf8;
            9'd203 : rom_q=8'h0;
            9'd204 : rom_q=8'hf8;
            9'd205 : rom_q=8'h0;
            9'd206 : rom_q=8'hf8;
            9'd207 : rom_q=8'h0;
            9'd208 : rom_q=8'hf8;
            9'd209 : rom_q=8'h0;
            9'd210 : rom_q=8'hf8;
            9'd211 : rom_q=8'h0;
            9'd212 : rom_q=8'hf8;
            9'd213 : rom_q=8'h0;
            9'd214 : rom_q=8'hf8;
            9'd215 : rom_q=8'h0;
            9'd216 : rom_q=8'hf8;
            9'd217 : rom_q=8'h0;
            9'd218 : rom_q=8'hf8;
            9'd219 : rom_q=8'h0;
            9'd220 : rom_q=8'hf8;
            9'd221 : rom_q=8'h0;
            9'd222 : rom_q=8'hf8;
            9'd223 : rom_q=8'h0;
            9'd224 : rom_q=8'hf8;
            9'd225 : rom_q=8'h0;
            9'd226 : rom_q=8'hf8;
            9'd227 : rom_q=8'h0;
            9'd228 : rom_q=8'hf8;
            9'd229 : rom_q=8'h0;
            9'd230 : rom_q=8'hf8;
            9'd231 : rom_q=8'h0;
            9'd232 : rom_q=8'hf8;
            9'd233 : rom_q=8'h0;
            9'd234 : rom_q=8'hf8;
            9'd235 : rom_q=8'h0;
            9'd236 : rom_q=8'hf8;
            9'd237 : rom_q=8'h0;
            9'd238 : rom_q=8'hf8;
            9'd239 : rom_q=8'h0;
            9'd240 : rom_q=8'h0;
            9'd241 : rom_q=8'h1F;
            9'd242 : rom_q=8'h0;
            9'd243 : rom_q=8'h1F;
            9'd244 : rom_q=8'h0;
            9'd245 : rom_q=8'h1F;
            9'd246 : rom_q=8'h0;
            9'd247 : rom_q=8'h1F;
            9'd248 : rom_q=8'h0;
            9'd249 : rom_q=8'h1F;
            9'd250 : rom_q=8'h0;
            9'd251 : rom_q=8'h1F;
            9'd252 : rom_q=8'h0;
            9'd253 : rom_q=8'h1F;
            9'd254 : rom_q=8'h0;
            9'd255 : rom_q=8'h1F;
            9'd256 : rom_q=8'h0;
            9'd257 : rom_q=8'h1F;
            9'd258 : rom_q=8'h0;
            9'd259 : rom_q=8'h1F;
            9'd260 : rom_q=8'h0;
            9'd261 : rom_q=8'h1F;
            9'd262 : rom_q=8'h0;
            9'd263 : rom_q=8'h1F;
            9'd264 : rom_q=8'h0;
            9'd265 : rom_q=8'h1F;
            9'd266 : rom_q=8'h0;
            9'd267 : rom_q=8'h1F;
            9'd268 : rom_q=8'h0;
            9'd269 : rom_q=8'h1F;
            9'd270 : rom_q=8'h0;
            9'd271 : rom_q=8'h1F;
            9'd272 : rom_q=8'h0;
            9'd273 : rom_q=8'h1F;
            9'd274 : rom_q=8'h0;
            9'd275 : rom_q=8'h1F;
            9'd276 : rom_q=8'h0;
            9'd277 : rom_q=8'h1F;
            9'd278 : rom_q=8'h0;
            9'd279 : rom_q=8'h1F;
            9'd280 : rom_q=8'h0;
            9'd281 : rom_q=8'h1F;
            9'd282 : rom_q=8'h0;
            9'd283 : rom_q=8'h1F;
            9'd284 : rom_q=8'h0;
            9'd285 : rom_q=8'h1F;
            9'd286 : rom_q=8'h0;
            9'd287 : rom_q=8'h1F;
            9'd288 : rom_q=8'h0;
            9'd289 : rom_q=8'h1F;
            9'd290 : rom_q=8'h0;
            9'd291 : rom_q=8'h1F;
            9'd292 : rom_q=8'h0;
            9'd293 : rom_q=8'h1F;
            9'd294 : rom_q=8'h0;
            9'd295 : rom_q=8'h1F;
            9'd296 : rom_q=8'h0;
            9'd297 : rom_q=8'h1F;
            9'd298 : rom_q=8'h0;
            9'd299 : rom_q=8'h1F;
            9'd300 : rom_q=8'h0;
            9'd301 : rom_q=8'h1F;
            9'd302 : rom_q=8'h0;
            9'd303 : rom_q=8'h1F;
            9'd304 : rom_q=8'h0;
            9'd305 : rom_q=8'h1F;
            9'd306 : rom_q=8'h0;
            9'd307 : rom_q=8'h1F;
            9'd308 : rom_q=8'h0;
            9'd309 : rom_q=8'h1F;
            9'd310 : rom_q=8'h0;
            9'd311 : rom_q=8'h1F;
            9'd312 : rom_q=8'h0;
            9'd313 : rom_q=8'h1F;
            9'd314 : rom_q=8'h0;
            9'd315 : rom_q=8'h1F;
            9'd316 : rom_q=8'h0;
            9'd317 : rom_q=8'h1F;
            9'd318 : rom_q=8'h0;
            9'd319 : rom_q=8'h1F;
            9'd320 : rom_q=8'h0;
            9'd321 : rom_q=8'h1F;
            9'd322 : rom_q=8'h0;
            9'd323 : rom_q=8'h1F;
            9'd324 : rom_q=8'h0;
            9'd325 : rom_q=8'h1F;
            9'd326 : rom_q=8'h0;
            9'd327 : rom_q=8'h1F;
            9'd328 : rom_q=8'h0;
            9'd329 : rom_q=8'h1F;
            9'd330 : rom_q=8'h0;
            9'd331 : rom_q=8'h1F;
            9'd332 : rom_q=8'h0;
            9'd333 : rom_q=8'h1F;
            9'd334 : rom_q=8'h0;
            9'd335 : rom_q=8'h1F;
            9'd336 : rom_q=8'h0;
            9'd337 : rom_q=8'h1F;
            9'd338 : rom_q=8'h0;
            9'd339 : rom_q=8'h1F;
            9'd340 : rom_q=8'h0;
            9'd341 : rom_q=8'h1F;
            9'd342 : rom_q=8'h0;
            9'd343 : rom_q=8'h1F;
            9'd344 : rom_q=8'h0;
            9'd345 : rom_q=8'h1F;
            9'd346 : rom_q=8'h0;
            9'd347 : rom_q=8'h1F;
            9'd348 : rom_q=8'h0;
            9'd349 : rom_q=8'h1F;
            9'd350 : rom_q=8'h0;
            9'd351 : rom_q=8'h1F;
            9'd352 : rom_q=8'h0;
            9'd353 : rom_q=8'h1F;
            9'd354 : rom_q=8'h0;
            9'd355 : rom_q=8'h1F;
            9'd356 : rom_q=8'h0;
            9'd357 : rom_q=8'h1F;
            9'd358 : rom_q=8'h0;
            9'd359 : rom_q=8'h1F;
            9'd360 : rom_q=8'h0;
            9'd361 : rom_q=8'h1F;
            9'd362 : rom_q=8'h0;
            9'd363 : rom_q=8'h1F;
            9'd364 : rom_q=8'h0;
            9'd365 : rom_q=8'h1F;
            9'd366 : rom_q=8'h0;
            9'd367 : rom_q=8'h1F;
            9'd368 : rom_q=8'h0;
            9'd369 : rom_q=8'h1F;
            9'd370 : rom_q=8'h0;
            9'd371 : rom_q=8'h1F;
            9'd372 : rom_q=8'h0;
            9'd373 : rom_q=8'h1F;
            9'd374 : rom_q=8'h0;
            9'd375 : rom_q=8'h1F;
            9'd376 : rom_q=8'h0;
            9'd377 : rom_q=8'h1F;
            9'd378 : rom_q=8'h0;
            9'd379 : rom_q=8'h1F;
            9'd380 : rom_q=8'h0;
            9'd381 : rom_q=8'h1F;
            9'd382 : rom_q=8'h0;
            9'd383 : rom_q=8'h1F;
            9'd384 : rom_q=8'h0;
            9'd385 : rom_q=8'h1F;
            9'd386 : rom_q=8'h0;
            9'd387 : rom_q=8'h1F;
            9'd388 : rom_q=8'h0;
            9'd389 : rom_q=8'h1F;
            9'd390 : rom_q=8'h0;
            9'd391 : rom_q=8'h1F;
            9'd392 : rom_q=8'h0;
            9'd393 : rom_q=8'h1F;
            9'd394 : rom_q=8'h0;
            9'd395 : rom_q=8'h1F;
            9'd396 : rom_q=8'h0;
            9'd397 : rom_q=8'h1F;
            9'd398 : rom_q=8'h0;
            9'd399 : rom_q=8'h1F;
            9'd400 : rom_q=8'h0;
            9'd401 : rom_q=8'h1F;
            9'd402 : rom_q=8'h0;
            9'd403 : rom_q=8'h1F;
            9'd404 : rom_q=8'h0;
            9'd405 : rom_q=8'h1F;
            9'd406 : rom_q=8'h0;
            9'd407 : rom_q=8'h1F;
            9'd408 : rom_q=8'h0;
            9'd409 : rom_q=8'h1F;
            9'd410 : rom_q=8'h0;
            9'd411 : rom_q=8'h1F;
            9'd412 : rom_q=8'h0;
            9'd413 : rom_q=8'h1F;
            9'd414 : rom_q=8'h0;
            9'd415 : rom_q=8'h1F;
            9'd416 : rom_q=8'h0;
            9'd417 : rom_q=8'h1F;
            9'd418 : rom_q=8'h0;
            9'd419 : rom_q=8'h1F;
            9'd420 : rom_q=8'h0;
            9'd421 : rom_q=8'h1F;
            9'd422 : rom_q=8'h0;
            9'd423 : rom_q=8'h1F;
            9'd424 : rom_q=8'h0;
            9'd425 : rom_q=8'h1F;
            9'd426 : rom_q=8'h0;
            9'd427 : rom_q=8'h1F;
            9'd428 : rom_q=8'h0;
            9'd429 : rom_q=8'h1F;
            9'd430 : rom_q=8'h0;
            9'd431 : rom_q=8'h1F;
            9'd432 : rom_q=8'h0;
            9'd433 : rom_q=8'h1F;
            9'd434 : rom_q=8'h0;
            9'd435 : rom_q=8'h1F;
            9'd436 : rom_q=8'h0;
            9'd437 : rom_q=8'h1F;
            9'd438 : rom_q=8'h0;
            9'd439 : rom_q=8'h1F;
            9'd440 : rom_q=8'h0;
            9'd441 : rom_q=8'h1F;
            9'd442 : rom_q=8'h0;
            9'd443 : rom_q=8'h1F;
            9'd444 : rom_q=8'h0;
            9'd445 : rom_q=8'h1F;
            9'd446 : rom_q=8'h0;
            9'd447 : rom_q=8'h1F;
            9'd448 : rom_q=8'h0;
            9'd449 : rom_q=8'h1F;
            9'd450 : rom_q=8'h0;
            9'd451 : rom_q=8'h1F;
            9'd452 : rom_q=8'h0;
            9'd453 : rom_q=8'h1F;
            9'd454 : rom_q=8'h0;
            9'd455 : rom_q=8'h1F;
            9'd456 : rom_q=8'h0;
            9'd457 : rom_q=8'h1F;
            9'd458 : rom_q=8'h0;
            9'd459 : rom_q=8'h1F;
            9'd460 : rom_q=8'h0;
            9'd461 : rom_q=8'h1F;
            9'd462 : rom_q=8'h0;
            9'd463 : rom_q=8'h1F;
            9'd464 : rom_q=8'h0;
            9'd465 : rom_q=8'h1F;
            9'd466 : rom_q=8'h0;
            9'd467 : rom_q=8'h1F;
            9'd468 : rom_q=8'h0;
            9'd469 : rom_q=8'h1F;
            9'd470 : rom_q=8'h0;
            9'd471 : rom_q=8'h1F;
            9'd472 : rom_q=8'h0;
            9'd473 : rom_q=8'h1F;
            9'd474 : rom_q=8'h0;
            9'd475 : rom_q=8'h1F;
            9'd476 : rom_q=8'h0;
            9'd477 : rom_q=8'h1F;
            9'd478 : rom_q=8'h0;
            9'd479 : rom_q=8'h1F;

            default: rom_q=8'd0;  
				
		endcase

endmodule
