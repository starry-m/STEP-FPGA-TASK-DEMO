
`timescale 1 ns / 100 ps
module pic_ram (address, q);

    input wire [8:0] address;
    output reg [239:0] q;
	 
	always @ (*)
		case(address)
			9'd0  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd1  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd2  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd3  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd4  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd5  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd6  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd7  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd8  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd9  : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd10 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd11 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd12 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd13 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd14 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd15 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd16 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd17 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd18 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd19 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd20 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd21 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd22 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd23 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd24 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd25 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd26 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd27 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd28 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd29 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd30 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd31 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd32 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd33 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd34 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd35 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd36 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd37 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd38 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd39 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd40 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd41 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd42 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd43 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd44 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd45 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd46 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd47 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd48 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd49 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd50 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd51 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd52 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd53 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd54 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd55 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd56 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd57 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd58 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd59 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd60 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd61 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd62 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd63 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd64 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd65 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd66 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd67 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd68 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd69 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd70 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd71 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd72 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd73 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd74 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd75 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd76 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd77 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd78 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd79 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd80 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd81 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd82 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd83 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd84 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd85 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd86 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd87 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd88 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd89 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd90 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd91 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd92 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd93 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd94 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd95 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd96 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd97 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd98 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd99 : q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd100: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd101: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd102: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd103: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd104: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd105: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd106: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd107: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd108: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd109: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd110: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd111: q = 240'h00000000000000000000000000000FF8000000000000000000000000000;
			9'd112: q = 240'h00000000000000000000000000003FFE000000000000000000000000000;
			9'd113: q = 240'h0000000000000000000000000000FFFF800000000000000000000000000;
			9'd114: q = 240'h0000000000000000000000000001FFFFC00000000000000000000000000;
			9'd115: q = 240'h0000000000000000000000000003FFFFE00000000000000000000000000;
			9'd116: q = 240'h0000000000000000000000000007FFFFF00000000000000000000000000;
			9'd117: q = 240'h000000000000000000000000000FFFFFF80000000000000000000000000;
			9'd118: q = 240'h000000000000000000000000000FFFFFF80000000000000000000000000;
			9'd119: q = 240'h000000000000000000000000001FFFFFFC0000000000000000000000000;
			9'd120: q = 240'h000000000000000000000000001FFFFFFC0000000000000000000000000;
			9'd121: q = 240'h000000000000000000000000001FFC1FFC0000000000000000000000000;
			9'd122: q = 240'h000000000000000000000000001FF80FFC0000000000000000000000000;
			9'd123: q = 240'h000000000000000000000000001FF00FFC0000000000000000000000000;
			9'd124: q = 240'h000000000000000000000000001FF007FC0000000000000000000000000;
			9'd125: q = 240'h000000000000000000000000001FF00FFC0000000000000000000000000;
			9'd126: q = 240'h000000000000000000000000001FF80FFC0000000000000000000000000;
			9'd127: q = 240'h000000000000000000000000001FF81FFC0000000000000000000000000;
			9'd128: q = 240'h000000000000000000000000001FFE3FFC0000000000000000000000000;
			9'd129: q = 240'h000000000000000000000000001FFE7FFC0000000000000000000000000;
			9'd130: q = 240'h000000000000000000000000000FFE7FF80000000000000000000000000;
			9'd131: q = 240'h000000000000000000000000000FFE7FF80000007FC0000000000000000;
			9'd132: q = 240'h0000000000000000000000000007FE7FF0000001FFF0000000000000000;
			9'd133: q = 240'h0000000000000000000380000007FE7FE0000007FFF8000000000000000;
			9'd134: q = 240'h0000000000000000001FF8000003FE7FC000000FFFFC000000000000000;
			9'd135: q = 240'h0000000000000000007FFE000003FE7FC000001FFFFE000000000000000;
			9'd136: q = 240'h000000000000000000FFFF000003FE7F8000003FFFFF000000000000000;
			9'd137: q = 240'h000000000000000001FFFF800001FC7F8000003FFFFF000000000000000;
			9'd138: q = 240'h000000000000000003FFFFC00001FC7F0000007FFFFF800000000000000;
			9'd139: q = 240'h000000000000000003FFFFC00000FC7F0000007FFBFF800000000000000;
			9'd140: q = 240'h000000000000000007FFFFE00000FCFF0000007FE0FFC00000000000000;
			9'd141: q = 240'h000000000000000007F83FE00000FCFE000000FFC07FC00000000000000;
			9'd142: q = 240'h00000000000000000FF01FE000007CFE000000FFC03FC00000000000000;
			9'd143: q = 240'h00000000000000000FF00FE000007CFE000000FFC03FC00000000000000;
			9'd144: q = 240'h00000000000000000FF00FE000007CFC000000FFC03FC00000000000000;
			9'd145: q = 240'h00000000000000000FF00FE000007CFC000000FFC07FC00000000000000;
			9'd146: q = 240'h00000000000000000FF01FE000007CFC000000FFC0FFC00000000000000;
			9'd147: q = 240'h000000000000000007F81FE000007CFC000001FF81FF800000000000000;
			9'd148: q = 240'h000000000000000007FE1FE000007CF8000001FF8FFF800000000000000;
			9'd149: q = 240'h000000000000000007FF1FE0000078F8000001FF1FFF000000000000000;
			9'd150: q = 240'h000000000000000003FF8FE0000078F8000001FE3FFF000000000000000;
			9'd151: q = 240'h000000000000000003FF8FE0000078F8000003FC7FFE000000000000000;
			9'd152: q = 240'h000000000000000001FFCFE0000079F8000003FCFFFC000000000000000;
			9'd153: q = 240'h000000000000000000FFC7E0000079F0000003F8FFF8000000000000000;
			9'd154: q = 240'h0000000000000000007FE7F0000079F0000007F1FFF0000000000000000;
			9'd155: q = 240'h0000000000000000001FE3F0000079F0000007E3FFE0000000000000000;
			9'd156: q = 240'h0000000000000000000FF3F0000079F000000FC7FFC0000000000000000;
			9'd157: q = 240'h00000000000000000003F1F0000071F000000FCFFF80000000000000000;
			9'd158: q = 240'h00000000000000000001F9F0000071F000001F8FFE00000000000000000;
			9'd159: q = 240'h00000000000000000000F8F0000071F000001F1FFC00000000000000000;
			9'd160: q = 240'h000000000000000000007CF0000071F000003E3FF800000000000000000;
			9'd161: q = 240'h000000000000000000003C780000F3F000003C7FE000000000000000000;
			9'd162: q = 240'h000000000000000000001E780000F3F0000078FFC000000000000000000;
			9'd163: q = 240'h000000000000000000001E380000F3F80000F8FF0000000000000000000;
			9'd164: q = 240'h000000000000000000000F3C0000F3F80000F1FE0000000000000000000;
			9'd165: q = 240'h00000000000000000000071C0001E3FC0001E3FC0000000000000000000;
			9'd166: q = 240'h00000000000000000000079C0003E3FC0003C7F80000000000000000000;
			9'd167: q = 240'h00000000000000000000038E0003E3FE00078FF00000000000000000000;
			9'd168: q = 240'h0000000000000000000003CF0007E1FF001F0FC00000000000000000000;
			9'd169: q = 240'h0000000000000000000001C7C00FE1FFC07F1F800000000000000000000;
			9'd170: q = 240'h0000000000000000000001E3E03FC1FFFFFE3F000000000000000000000;
			9'd171: q = 240'h0000000000000000000000F3FFFFC8FFFFFC7E000000000000000000000;
			9'd172: q = 240'h0000000000000000000000F1FFFF8CFFFFF0FC000000000000000000000;
			9'd173: q = 240'h0000000000000000000000F8FFFF1C7FFFE1FC000000000000000000000;
			9'd174: q = 240'h00000000000000000000007C3FFE1E3FFFC3F8000000000000000000000;
			9'd175: q = 240'h00000000000000000000007E1FF83F1FFF07F0000000000000000000000;
			9'd176: q = 240'h00000000000000000000003F0000FF83FC0FE0000000000000000000000;
			9'd177: q = 240'h00000000000000000000003FC003FFC0003FC0000000000000000000000;
			9'd178: q = 240'h00000000000000000000001FF00FFFF000FFC0000000000000000000000;
			9'd179: q = 240'h00000000000000000000001FFFFFFFFE07FF80000000000000000000000;
			9'd180: q = 240'h00000000000000000000000FFFFFFFFFFFFF80000000000000000000000;
			9'd181: q = 240'h00000000000000000000000FFFFFFFFFFFFF00000000000000000000000;
			9'd182: q = 240'h000000000000000000000007FFFFFFFFFFFE00000000000000000000000;
			9'd183: q = 240'h000000000000000000000007FFFFFFFFFFFE00000000000000000000000;
			9'd184: q = 240'h000000000000000000000007FFFFFFFFFFFC00000000000000000000000;
			9'd185: q = 240'h000000000000000000000003FFFFFFFFFFFC00000000000000000000000;
			9'd186: q = 240'h000000000000000000000003FFFFFFFFFFFC00000000000000000000000;
			9'd187: q = 240'h000000000000000000000003FFFFFFFFFFF800000000000000000000000;
			9'd188: q = 240'h000000000000000000000001FFFFFFFFFFF800000000000000000000000;
			9'd189: q = 240'h000000000000000000000001FFFFFFFFFFF000000000000000000000000;
			9'd190: q = 240'h000000000000000000000000FFFFFFFFFFF000000000000000000000000;
			9'd191: q = 240'h000000000000000000000000FFFFFFFFFFF000000000000000000000000;
			9'd192: q = 240'h000000000000000000000000FFFFFFFFFFE000000000000000000000000;
			9'd193: q = 240'h0000000000000000000000007FFFFFFFFFE000000000000000000000000;
			9'd194: q = 240'h0000000000000000000000007FFFFFFFFFC000000000000000000000000;
			9'd195: q = 240'h0000000000000000000000007FFFFFFFFFC000000000000000000000000;
			9'd196: q = 240'h0000000000000000000000003FFFFFFFFFC000000000000000000000000;
			9'd197: q = 240'h0000000000000000000000003FFFFFFFFF8000000000000000000000000;
			9'd198: q = 240'h0000000000000000000000003FFFFFFFFF8000000000000000000000000;
			9'd199: q = 240'h0000000000000000000000001FFFFFFFFF8000000000000000000000000;
			9'd200: q = 240'h0000000000000000000000001FFFFFFFFF0000000000000000000000000;
			9'd201: q = 240'h0000000000000000000000001FFFFFFFFF0000000000000000000000000;
			9'd202: q = 240'h0000000000000000000000000FFFFFFFFE0000000000000000000000000;
			9'd203: q = 240'h0000000000000000000000000FFFFFFFFE0000000000000000000000000;
			9'd204: q = 240'h00000000000000000000000007FFFFFFFC0000000000000000000000000;
			9'd205: q = 240'h00000000000000000000000003FFFFFFFC0000000000000000000000000;
			9'd206: q = 240'h00000000000000000000000003FFFFFFF80000000000000000000000000;
			9'd207: q = 240'h00000000000000000000000001FFFFFFF00000000000000000000000000;
			9'd208: q = 240'h00000000000000000000000000FFFFFFE00000000000000000000000000;
			9'd209: q = 240'h000000000000000000000000007FFFFFC00000000000000000000000000;
			9'd210: q = 240'h000000000000000000000000003FFFFF800000000000000000000000000;
			9'd211: q = 240'h000000000000000000000000000FFFFE000000000000000000000000000;
			9'd212: q = 240'h0000000000000000000000000001FFF8000000000000000000000000000;
			9'd213: q = 240'h00000000000000000000000000003F80000000000000000000000000000;
			9'd214: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd215: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd216: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd217: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd218: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd219: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd220: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd221: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd222: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd223: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd224: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd225: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd226: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd227: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd228: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd229: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd230: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd231: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd232: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd233: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd234: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd235: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd236: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd237: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd238: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd239: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd230: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd241: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd242: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd243: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd244: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd245: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd246: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd247: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd248: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd249: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd250: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd251: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd252: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd253: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd254: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd255: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd256: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd257: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd258: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd259: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd260: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd261: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd262: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd263: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd264: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd265: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd266: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd267: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd268: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd269: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd270: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd271: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd272: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd273: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd274: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd275: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd276: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd277: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd278: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd279: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd280: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd281: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd282: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd283: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd284: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd285: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd286: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd287: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd288: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd289: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd290: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd291: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd292: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd293: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd294: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd295: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd296: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd297: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd298: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd299: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd300: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd301: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd302: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd303: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd304: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd305: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd306: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd307: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd308: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd309: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd310: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd311: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd312: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd313: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd314: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd315: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd316: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd317: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd318: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			9'd319: q = 240'h00000000000000000000000000000000000000000000000000000000000;
			default:q = 0;
			
			
			
		endcase
		
endmodule
