`timescale 1 ns / 100 ps
module lcd_ram(
        output reg [7:0] rom_q,
        input wire [8:0] rom_addr
);
	always @ (*)
		case(rom_addr)
            9'd0 : rom_q=8'd2;
            9'd1 : rom_q=8'd1;
            9'd2 : rom_q=8'd2;
            9'd3 : rom_q=8'd3;
            9'd4 : rom_q=8'd4;
            9'd5 : rom_q=8'd5;
            9'd6 : rom_q=8'd6;
            9'd7 : rom_q=8'd7;
            9'd8 : rom_q=8'd8;
            9'd9 : rom_q=8'd9;
            9'd10 : rom_q=8'd10;
            9'd11 : rom_q=8'd11;
            9'd12 : rom_q=8'd12;
            9'd13 : rom_q=8'd13;
            9'd14 : rom_q=8'd14;
            9'd15 : rom_q=8'd15;
            9'd16 : rom_q=8'd16;
            9'd17 : rom_q=8'd17;
            9'd18 : rom_q=8'd18;
            9'd19 : rom_q=8'd19;
            9'd20 : rom_q=8'd20;
            9'd21 : rom_q=8'd21;
            9'd22 : rom_q=8'd22;
            9'd23 : rom_q=8'd23;
            9'd24 : rom_q=8'd24;
            9'd25 : rom_q=8'd25;
            9'd26 : rom_q=8'd26;
            9'd27 : rom_q=8'd27;
            9'd28 : rom_q=8'd28;
            9'd29 : rom_q=8'd29;
            9'd30 : rom_q=8'd30;
            9'd31 : rom_q=8'd31;
            9'd32 : rom_q=8'd32;
            9'd33 : rom_q=8'd33;
            9'd34 : rom_q=8'd34;
            9'd35 : rom_q=8'd35;
            9'd36 : rom_q=8'd36;
            9'd37 : rom_q=8'd37;
            9'd38 : rom_q=8'd38;
            9'd39 : rom_q=8'd39;
            9'd40 : rom_q=8'd40;
            9'd41 : rom_q=8'd41;
            9'd42 : rom_q=8'd42;
            9'd43 : rom_q=8'd43;
            9'd44 : rom_q=8'd44;
            9'd45 : rom_q=8'd45;
            9'd46 : rom_q=8'd46;
            9'd47 : rom_q=8'd47;
            9'd48 : rom_q=8'd48;
            9'd49 : rom_q=8'd49;
            9'd50 : rom_q=8'd50;
            9'd51 : rom_q=8'd51;
            9'd52 : rom_q=8'd52;
            9'd53 : rom_q=8'd53;
            9'd54 : rom_q=8'd54;
            9'd55 : rom_q=8'd55;
            9'd56 : rom_q=8'd56;
            9'd57 : rom_q=8'd57;
            9'd58 : rom_q=8'd58;
            9'd59 : rom_q=8'd59;
            9'd60 : rom_q=8'd60;
            9'd61 : rom_q=8'd61;
            9'd62 : rom_q=8'd62;
            9'd63 : rom_q=8'd63;
            9'd64 : rom_q=8'd64;
            9'd65 : rom_q=8'd65;
            9'd66 : rom_q=8'd66;
            9'd67 : rom_q=8'd67;
            9'd68 : rom_q=8'd68;
            9'd69 : rom_q=8'd69;
            9'd70 : rom_q=8'd70;
            9'd71 : rom_q=8'd71;
            9'd72 : rom_q=8'd72;
            9'd73 : rom_q=8'd73;
            9'd74 : rom_q=8'd74;
            9'd75 : rom_q=8'd75;
            9'd76 : rom_q=8'd76;
            9'd77 : rom_q=8'd77;
            9'd78 : rom_q=8'd78;
            9'd79 : rom_q=8'd79;
            9'd80 : rom_q=8'd80;
            9'd81 : rom_q=8'd81;
            9'd82 : rom_q=8'd82;
            9'd83 : rom_q=8'd83;
            9'd84 : rom_q=8'd84;
            9'd85 : rom_q=8'd85;
            9'd86 : rom_q=8'd86;
            9'd87 : rom_q=8'd87;
            9'd88 : rom_q=8'd88;
            9'd89 : rom_q=8'd89;
            9'd90 : rom_q=8'd90;
            9'd91 : rom_q=8'd91;
            9'd92 : rom_q=8'd92;
            9'd93 : rom_q=8'd93;
            9'd94 : rom_q=8'd94;
            9'd95 : rom_q=8'd95;
            9'd96 : rom_q=8'd96;
            9'd97 : rom_q=8'd97;
            9'd98 : rom_q=8'd98;
            9'd99 : rom_q=8'd99;
            9'd100 : rom_q=8'd100;
            9'd101 : rom_q=8'd101;
            9'd102 : rom_q=8'd102;
            9'd103 : rom_q=8'd103;
            9'd104 : rom_q=8'd104;
            9'd105 : rom_q=8'd105;
            9'd106 : rom_q=8'd106;
            9'd107 : rom_q=8'd107;
            9'd108 : rom_q=8'd108;
            9'd109 : rom_q=8'd109;
            9'd110 : rom_q=8'd110;
            9'd111 : rom_q=8'd111;
            9'd112 : rom_q=8'd112;
            9'd113 : rom_q=8'd113;
            9'd114 : rom_q=8'd114;
            9'd115 : rom_q=8'd115;
            9'd116 : rom_q=8'd116;
            9'd117 : rom_q=8'd117;
            9'd118 : rom_q=8'd118;
            9'd119 : rom_q=8'd119;
            9'd120 : rom_q=8'd120;
            9'd121 : rom_q=8'd121;
            9'd122 : rom_q=8'd122;
            9'd123 : rom_q=8'd123;
            9'd124 : rom_q=8'd124;
            9'd125 : rom_q=8'd125;
            9'd126 : rom_q=8'd126;
            9'd127 : rom_q=8'd127;
            9'd128 : rom_q=8'd128;
            9'd129 : rom_q=8'd129;
            9'd130 : rom_q=8'd130;
            9'd131 : rom_q=8'd131;
            9'd132 : rom_q=8'd132;
            9'd133 : rom_q=8'd133;
            9'd134 : rom_q=8'd134;
            9'd135 : rom_q=8'd135;
            9'd136 : rom_q=8'd136;
            9'd137 : rom_q=8'd137;
            9'd138 : rom_q=8'd138;
            9'd139 : rom_q=8'd139;
            9'd140 : rom_q=8'd140;
            9'd141 : rom_q=8'd141;
            9'd142 : rom_q=8'd142;
            9'd143 : rom_q=8'd143;
            9'd144 : rom_q=8'd144;
            9'd145 : rom_q=8'd145;
            9'd146 : rom_q=8'd146;
            9'd147 : rom_q=8'd147;
            9'd148 : rom_q=8'd148;
            9'd149 : rom_q=8'd149;
            9'd150 : rom_q=8'd150;
            9'd151 : rom_q=8'd151;
            9'd152 : rom_q=8'd152;
            9'd153 : rom_q=8'd153;
            9'd154 : rom_q=8'd154;
            9'd155 : rom_q=8'd155;
            9'd156 : rom_q=8'd156;
            9'd157 : rom_q=8'd157;
            9'd158 : rom_q=8'd158;
            9'd159 : rom_q=8'd159;
            9'd160 : rom_q=8'd160;
            9'd161 : rom_q=8'd161;
            9'd162 : rom_q=8'd162;
            9'd163 : rom_q=8'd163;
            9'd164 : rom_q=8'd164;
            9'd165 : rom_q=8'd165;
            9'd166 : rom_q=8'd166;
            9'd167 : rom_q=8'd167;
            9'd168 : rom_q=8'd168;
            9'd169 : rom_q=8'd169;
            9'd170 : rom_q=8'd170;
            9'd171 : rom_q=8'd171;
            9'd172 : rom_q=8'd172;
            9'd173 : rom_q=8'd173;
            9'd174 : rom_q=8'd174;
            9'd175 : rom_q=8'd175;
            9'd176 : rom_q=8'd176;
            9'd177 : rom_q=8'd177;
            9'd178 : rom_q=8'd178;
            9'd179 : rom_q=8'd179;
            9'd180 : rom_q=8'd180;
            9'd181 : rom_q=8'd181;
            9'd182 : rom_q=8'd182;
            9'd183 : rom_q=8'd183;
            9'd184 : rom_q=8'd184;
            9'd185 : rom_q=8'd185;
            9'd186 : rom_q=8'd186;
            9'd187 : rom_q=8'd187;
            9'd188 : rom_q=8'd188;
            9'd189 : rom_q=8'd189;
            9'd190 : rom_q=8'd190;
            9'd191 : rom_q=8'd191;
            9'd192 : rom_q=8'd192;
            9'd193 : rom_q=8'd193;
            9'd194 : rom_q=8'd194;
            9'd195 : rom_q=8'd195;
            9'd196 : rom_q=8'd196;
            9'd197 : rom_q=8'd197;
            9'd198 : rom_q=8'd198;
            9'd199 : rom_q=8'd199;
            9'd200 : rom_q=8'd200;
            9'd201 : rom_q=8'd201;
            9'd202 : rom_q=8'd202;
            9'd203 : rom_q=8'd203;
            9'd204 : rom_q=8'd204;
            9'd205 : rom_q=8'd205;
            9'd206 : rom_q=8'd206;
            9'd207 : rom_q=8'd207;
            9'd208 : rom_q=8'd208;
            9'd209 : rom_q=8'd209;
            9'd210 : rom_q=8'd210;
            9'd211 : rom_q=8'd211;
            9'd212 : rom_q=8'd212;
            9'd213 : rom_q=8'd213;
            9'd214 : rom_q=8'd214;
            9'd215 : rom_q=8'd215;
            9'd216 : rom_q=8'd216;
            9'd217 : rom_q=8'd217;
            9'd218 : rom_q=8'd218;
            9'd219 : rom_q=8'd219;
            9'd220 : rom_q=8'd220;
            9'd221 : rom_q=8'd221;
            9'd222 : rom_q=8'd222;
            9'd223 : rom_q=8'd223;
            9'd224 : rom_q=8'd224;
            9'd225 : rom_q=8'd225;
            9'd226 : rom_q=8'd226;
            9'd227 : rom_q=8'd227;
            9'd228 : rom_q=8'd228;
            9'd229 : rom_q=8'd229;
            9'd230 : rom_q=8'd230;
            9'd231 : rom_q=8'd231;
            9'd232 : rom_q=8'd232;
            9'd233 : rom_q=8'd233;
            9'd234 : rom_q=8'd234;
            9'd235 : rom_q=8'd235;
            9'd236 : rom_q=8'd236;
            9'd237 : rom_q=8'd237;
            9'd238 : rom_q=8'd238;
            9'd239 : rom_q=8'd239;
            9'd240 : rom_q=8'd240;
            9'd241 : rom_q=8'd241;
            9'd242 : rom_q=8'd242;
            9'd243 : rom_q=8'd243;
            9'd244 : rom_q=8'd244;
            9'd245 : rom_q=8'd245;
            9'd246 : rom_q=8'd246;
            9'd247 : rom_q=8'd247;
            9'd248 : rom_q=8'd248;
            9'd249 : rom_q=8'd249;
            9'd250 : rom_q=8'd250;
            9'd251 : rom_q=8'd251;
            9'd252 : rom_q=8'd252;
            9'd253 : rom_q=8'd253;
            9'd254 : rom_q=8'd254;
            9'd255 : rom_q=8'd255;
            9'd256 : rom_q=8'd0;
            9'd257 : rom_q=8'd1;
            9'd258 : rom_q=8'd2;
            9'd259 : rom_q=8'd3;
            9'd260 : rom_q=8'd4;
            9'd261 : rom_q=8'd5;
            9'd262 : rom_q=8'd6;
            9'd263 : rom_q=8'd7;
            9'd264 : rom_q=8'd8;
            9'd265 : rom_q=8'd9;
            9'd266 : rom_q=8'd10;
            9'd267 : rom_q=8'd11;
            9'd268 : rom_q=8'd12;
            9'd269 : rom_q=8'd13;
            9'd270 : rom_q=8'd14;
            9'd271 : rom_q=8'd15;
            9'd272 : rom_q=8'd16;
            9'd273 : rom_q=8'd17;
            9'd274 : rom_q=8'd18;
            9'd275 : rom_q=8'd19;
            9'd276 : rom_q=8'd20;
            9'd277 : rom_q=8'd21;
            9'd278 : rom_q=8'd22;
            9'd279 : rom_q=8'd23;
            9'd280 : rom_q=8'd24;
            9'd281 : rom_q=8'd25;
            9'd282 : rom_q=8'd26;
            9'd283 : rom_q=8'd27;
            9'd284 : rom_q=8'd28;
            9'd285 : rom_q=8'd29;
            9'd286 : rom_q=8'd30;
            9'd287 : rom_q=8'd31;
            9'd288 : rom_q=8'd32;
            9'd289 : rom_q=8'd33;
            9'd290 : rom_q=8'd34;
            9'd291 : rom_q=8'd35;
            9'd292 : rom_q=8'd36;
            9'd293 : rom_q=8'd37;
            9'd294 : rom_q=8'd38;
            9'd295 : rom_q=8'd39;
            9'd296 : rom_q=8'd40;
            9'd297 : rom_q=8'd41;
            9'd298 : rom_q=8'd42;
            9'd299 : rom_q=8'd43;
            9'd300 : rom_q=8'd44;
            9'd301 : rom_q=8'd45;
            9'd302 : rom_q=8'd46;
            9'd303 : rom_q=8'd47;
            9'd304 : rom_q=8'd48;
            9'd305 : rom_q=8'd49;
            9'd306 : rom_q=8'd50;
            9'd307 : rom_q=8'd51;
            9'd308 : rom_q=8'd52;
            9'd309 : rom_q=8'd53;
            9'd310 : rom_q=8'd54;
            9'd311 : rom_q=8'd55;
            9'd312 : rom_q=8'd56;
            9'd313 : rom_q=8'd57;
            9'd314 : rom_q=8'd58;
            9'd315 : rom_q=8'd59;
            9'd316 : rom_q=8'd60;
            9'd317 : rom_q=8'd61;
            9'd318 : rom_q=8'd62;
            9'd319 : rom_q=8'd63;
            9'd320 : rom_q=8'd64;
            9'd321 : rom_q=8'd65;
            9'd322 : rom_q=8'd66;
            9'd323 : rom_q=8'd67;
            9'd324 : rom_q=8'd68;
            9'd325 : rom_q=8'd69;
            9'd326 : rom_q=8'd70;
            9'd327 : rom_q=8'd71;
            9'd328 : rom_q=8'd72;
            9'd329 : rom_q=8'd73;
            9'd330 : rom_q=8'd74;
            9'd331 : rom_q=8'd75;
            9'd332 : rom_q=8'd76;
            9'd333 : rom_q=8'd77;
            9'd334 : rom_q=8'd78;
            9'd335 : rom_q=8'd79;
            9'd336 : rom_q=8'd80;
            9'd337 : rom_q=8'd81;
            9'd338 : rom_q=8'd82;
            9'd339 : rom_q=8'd83;
            9'd340 : rom_q=8'd84;
            9'd341 : rom_q=8'd85;
            9'd342 : rom_q=8'd86;
            9'd343 : rom_q=8'd87;
            9'd344 : rom_q=8'd88;
            9'd345 : rom_q=8'd89;
            9'd346 : rom_q=8'd90;
            9'd347 : rom_q=8'd91;
            9'd348 : rom_q=8'd92;
            9'd349 : rom_q=8'd93;
            9'd350 : rom_q=8'd94;
            9'd351 : rom_q=8'd95;
            9'd352 : rom_q=8'd96;
            9'd353 : rom_q=8'd97;
            9'd354 : rom_q=8'd98;
            9'd355 : rom_q=8'd99;
            9'd356 : rom_q=8'd100;
            9'd357 : rom_q=8'd101;
            9'd358 : rom_q=8'd102;
            9'd359 : rom_q=8'd103;
            9'd360 : rom_q=8'd104;
            9'd361 : rom_q=8'd105;
            9'd362 : rom_q=8'd106;
            9'd363 : rom_q=8'd107;
            9'd364 : rom_q=8'd108;
            9'd365 : rom_q=8'd109;
            9'd366 : rom_q=8'd110;
            9'd367 : rom_q=8'd111;
            9'd368 : rom_q=8'd112;
            9'd369 : rom_q=8'd113;
            9'd370 : rom_q=8'd114;
            9'd371 : rom_q=8'd115;
            9'd372 : rom_q=8'd116;
            9'd373 : rom_q=8'd117;
            9'd374 : rom_q=8'd118;
            9'd375 : rom_q=8'd119;
            9'd376 : rom_q=8'd120;
            9'd377 : rom_q=8'd121;
            9'd378 : rom_q=8'd122;
            9'd379 : rom_q=8'd123;
            9'd380 : rom_q=8'd124;
            9'd381 : rom_q=8'd125;
            9'd382 : rom_q=8'd126;
            9'd383 : rom_q=8'd127;
            9'd384 : rom_q=8'd128;
            9'd385 : rom_q=8'd129;
            9'd386 : rom_q=8'd130;
            9'd387 : rom_q=8'd131;
            9'd388 : rom_q=8'd132;
            9'd389 : rom_q=8'd133;
            9'd390 : rom_q=8'd134;
            9'd391 : rom_q=8'd135;
            9'd392 : rom_q=8'd136;
            9'd393 : rom_q=8'd137;
            9'd394 : rom_q=8'd138;
            9'd395 : rom_q=8'd139;
            9'd396 : rom_q=8'd140;
            9'd397 : rom_q=8'd141;
            9'd398 : rom_q=8'd142;
            9'd399 : rom_q=8'd143;
            9'd400 : rom_q=8'd144;
            9'd401 : rom_q=8'd145;
            9'd402 : rom_q=8'd146;
            9'd403 : rom_q=8'd147;
            9'd404 : rom_q=8'd148;
            9'd405 : rom_q=8'd149;
            9'd406 : rom_q=8'd150;
            9'd407 : rom_q=8'd151;
            9'd408 : rom_q=8'd152;
            9'd409 : rom_q=8'd153;
            9'd410 : rom_q=8'd154;
            9'd411 : rom_q=8'd155;
            9'd412 : rom_q=8'd156;
            9'd413 : rom_q=8'd157;
            9'd414 : rom_q=8'd158;
            9'd415 : rom_q=8'd159;
            9'd416 : rom_q=8'd160;
            9'd417 : rom_q=8'd161;
            9'd418 : rom_q=8'd162;
            9'd419 : rom_q=8'd163;
            9'd420 : rom_q=8'd164;
            9'd421 : rom_q=8'd165;
            9'd422 : rom_q=8'd166;
            9'd423 : rom_q=8'd167;
            9'd424 : rom_q=8'd168;
            9'd425 : rom_q=8'd169;
            9'd426 : rom_q=8'd170;
            9'd427 : rom_q=8'd171;
            9'd428 : rom_q=8'd172;
            9'd429 : rom_q=8'd173;
            9'd430 : rom_q=8'd174;
            9'd431 : rom_q=8'd175;
            9'd432 : rom_q=8'd176;
            9'd433 : rom_q=8'd177;
            9'd434 : rom_q=8'd178;
            9'd435 : rom_q=8'd179;
            9'd436 : rom_q=8'd180;
            9'd437 : rom_q=8'd181;
            9'd438 : rom_q=8'd182;
            9'd439 : rom_q=8'd183;
            9'd440 : rom_q=8'd184;
            9'd441 : rom_q=8'd185;
            9'd442 : rom_q=8'd186;
            9'd443 : rom_q=8'd187;
            9'd444 : rom_q=8'd188;
            9'd445 : rom_q=8'd189;
            9'd446 : rom_q=8'd190;
            9'd447 : rom_q=8'd191;
            9'd448 : rom_q=8'd192;
            9'd449 : rom_q=8'd193;
            9'd450 : rom_q=8'd194;
            9'd451 : rom_q=8'd195;
            9'd452 : rom_q=8'd196;
            9'd453 : rom_q=8'd197;
            9'd454 : rom_q=8'd198;
            9'd455 : rom_q=8'd199;
            9'd456 : rom_q=8'd200;
            9'd457 : rom_q=8'd201;
            9'd458 : rom_q=8'd202;
            9'd459 : rom_q=8'd203;
            9'd460 : rom_q=8'd204;
            9'd461 : rom_q=8'd205;
            9'd462 : rom_q=8'd206;
            9'd463 : rom_q=8'd207;
            9'd464 : rom_q=8'd208;
            9'd465 : rom_q=8'd209;
            9'd466 : rom_q=8'd210;
            9'd467 : rom_q=8'd211;
            9'd468 : rom_q=8'd212;
            9'd469 : rom_q=8'd213;
            9'd470 : rom_q=8'd214;
            9'd471 : rom_q=8'd215;
            9'd472 : rom_q=8'd216;
            9'd473 : rom_q=8'd217;
            9'd474 : rom_q=8'd218;
            9'd475 : rom_q=8'd219;
            9'd476 : rom_q=8'd220;
            9'd477 : rom_q=8'd221;
            9'd478 : rom_q=8'd222;
            9'd479 : rom_q=8'd223;   
            default: rom_q=8'd0;  
				
		endcase

endmodule
